//MODULOS
module GNOT(a,x);
	input a;
	output x;

//ASIGNACIONES
assign x=~a;
endmodule
