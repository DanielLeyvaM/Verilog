module Display(sw,a_to_g);
	input [3:0] sw;
	output [6:0] a_to_g;
	
assign a_to_g = 
		(sw==0)? 7'b100_0000:
		(sw==1)? 7'b111_1001:
		(sw==2)? 7'b010_0100:
		(sw==3)? 7'b011_0000:
		(sw==4)? 7'b001_1001:
		(sw==5)? 7'b001_0010:
		(sw==6)? 7'b000_0010:
		(sw==7)? 7'b111_1000:
		(sw==8)? 7'b000_0000:
		(sw==9)? 7'b001_0000:
		(sw=='hA)? 7'b000_1000:
		(sw=='hB)? 7'b000_0011:
		(sw=='hC)? 7'b100_0110:
		(sw=='hD)? 7'b010_0001:
		(sw=='hE)? 7'b000_0110:
		           7'b000_1110;
endmodule
